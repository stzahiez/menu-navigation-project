work.sync_rst_gen(rtl_sync_rst_gen) :[0[:
work.altsyncram(altsyncram) rtlc_no_parameters
work.general_fifo(arc_general_fifo) :[0[: :8: :640: :10: :8: :1:
work.debouncer(debouncer_rtl) :50000000: :[0[:
work.checksum_calc(arc_checksum_calc) :[0[: :false: :0: :8: :8:
work.ram_simple(arc_ram_simple) :[0[: :8: :10:
work.wbs_reg(rtl_wbs_reg) :[0[: :8: :4:
work.hexss(arc_hexss) rtlc_no_parameters
